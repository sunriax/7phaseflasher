.title KiCad schematic
R17 Net-_C3-Pad1_ GND 47k
D2 GND Net-_D2-Pad2_ LED
C2 Net-_C2-Pad1_ GND 10u
C3 Net-_C3-Pad1_ GND 10u
Q2 Net-_C2-Pad1_ Net-_Q2-Pad2_ Net-_D2-Pad2_ BC547
R9 Net-_Q2-Pad2_ Net-_C3-Pad1_ 47k
R2 +9V Net-_Q2-Pad2_ 470
C5 Net-_C5-Pad1_ GND 10u
R12 Net-_Q5-Pad2_ Net-_C6-Pad1_ 47k
C6 Net-_C6-Pad1_ GND 10u
R20 Net-_C6-Pad1_ GND 47k
Q5 Net-_C5-Pad1_ Net-_Q5-Pad2_ unconnected-_Q5-Pad3_ BC547
R5 +9V Net-_Q5-Pad2_ 470
R14 Net-_Q7-Pad2_ Net-_C1-Pad1_ 47k
R11 Net-_Q4-Pad2_ Net-_C5-Pad1_ 47k
R4 +9V Net-_Q4-Pad2_ 470
R19 Net-_C5-Pad1_ GND 47k
R18 Net-_C4-Pad1_ GND 47k
D3 GND Net-_D3-Pad2_ LED
Q3 Net-_C3-Pad1_ Net-_Q3-Pad2_ Net-_D3-Pad2_ BC547
D4 GND Net-_D4-Pad2_ LED
Q4 Net-_C4-Pad1_ Net-_Q4-Pad2_ Net-_D4-Pad2_ BC547
C4 Net-_C4-Pad1_ GND 10u
R3 +9V Net-_Q3-Pad2_ 470
R10 Net-_Q3-Pad2_ Net-_C4-Pad1_ 47k
R6 +9V Net-_Q6-Pad2_ 470
Q6 Net-_C6-Pad1_ Net-_Q6-Pad2_ Net-_D5-Pad2_ BC547
D6 GND Net-_D6-Pad2_ LED
C7 Net-_C7-Pad1_ GND 10u
R7 +9V Net-_Q7-Pad2_ 470
Q7 Net-_C7-Pad1_ Net-_Q7-Pad2_ Net-_D6-Pad2_ BC547
D5 GND Net-_D5-Pad2_ LED
R21 Net-_C7-Pad1_ GND 47k
R13 Net-_Q6-Pad2_ Net-_C7-Pad1_ 47k
R8 Net-_Q1-Pad2_ Net-_C2-Pad1_ 47k
C1 Net-_C1-Pad1_ GND 10u
R15 Net-_C1-Pad1_ GND 47k
Q1 Net-_C1-Pad1_ Net-_Q1-Pad2_ Net-_D1-Pad2_ BC547
J1 +9V Connector
R1 +9V Net-_Q1-Pad2_ 470
R16 Net-_C2-Pad1_ GND 47k
D1 GND Net-_D1-Pad2_ LED
J2 GND Connector
.end
